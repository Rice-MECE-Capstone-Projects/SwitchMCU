`timescale 1ns/1ps

module tb_smoke_riscv32i;

    // -----------------------------------------
    // Clock + GPIO
    // -----------------------------------------
    logic clk = 0;

    logic [31:0] GPIO0_R0_CH1;
    logic [31:0] GPIO0_R0_CH2;
    logic [31:0] GPIO0_R1_CH1;
    logic [31:0] GPIO0_R1_CH2;

    wire  STOP_sim;

    // -----------------------------------------
    // Data memory BRAM ports
    // -----------------------------------------
    wire        data_mem_clkb;
    wire        data_mem_enb;
    wire        data_mem_rstb;
    wire [3:0]  data_mem_web;
    wire [31:0] data_mem_addrb;
    wire [31:0] data_mem_dinb;
    wire        data_mem_rstb_busy;
    wire [31:0] data_mem_doutb;

    // -----------------------------------------
    // Instruction memory BRAM ports
    // -----------------------------------------
    wire        ins_mem_clkb;
    wire        ins_mem_enb;
    wire        ins_mem_rstb;
    wire [3:0]  ins_mem_web;
    wire [31:0] ins_mem_addrb;
    wire [31:0] ins_mem_dinb;
    wire        ins_mem_rstb_busy;
    wire [31:0] ins_mem_doutb;

    // -----------------------------------------
    // DUT
    // -----------------------------------------
    riscv32i dut (
        .clk(clk),

        .GPIO0_R0_CH1(GPIO0_R0_CH1),
        .GPIO0_R0_CH2(GPIO0_R0_CH2),
        .GPIO0_R1_CH1(GPIO0_R1_CH1),
        .GPIO0_R1_CH2(GPIO0_R1_CH2),
        .STOP_sim(STOP_sim),

        .data_mem_clkb(data_mem_clkb),
        .data_mem_enb(data_mem_enb),
        .data_mem_rstb(data_mem_rstb),
        .data_mem_web(data_mem_web),
        .data_mem_addrb(data_mem_addrb),
        .data_mem_dinb(data_mem_dinb),
        .data_mem_rstb_busy(data_mem_rstb_busy),
        .data_mem_doutb(data_mem_doutb),

        .ins_mem_clkb(ins_mem_clkb),
        .ins_mem_enb(ins_mem_enb),
        .ins_mem_rstb(ins_mem_rstb),
        .ins_mem_web(ins_mem_web),
        .ins_mem_addrb(ins_mem_addrb),
        .ins_mem_dinb(ins_mem_dinb),
        .ins_mem_rstb_busy(ins_mem_rstb_busy),
        .ins_mem_doutb(ins_mem_doutb)
    );

    // -----------------------------------------
    // Clock
    // -----------------------------------------
    always #5 clk = ~clk;


    // -----------------------------------------
    // Stimulus
    // -----------------------------------------
    initial begin
        $display("---- Smoke Test Start ----");

        GPIO0_R0_CH1 = 32'h0;
        GPIO0_R0_CH2 = 32'h00000600;
        GPIO0_R1_CH1 = 32'h00000384;
        GPIO0_R1_CH2 = 32'hDEADBEEF;

        repeat (10) @(posedge clk);

        // Reset pulse
        GPIO0_R0_CH1 = 32'b10;
        @(posedge clk);
        GPIO0_R0_CH1 = 32'b00;

        // Start pulse
        @(posedge clk);
        GPIO0_R0_CH1 = 32'b01;
        @(posedge clk);

        // Run until timeout
        repeat (2000) @(posedge clk);
        $display("TIMEOUT: Simulation stopped.");
        $finish;
    end

    // -------------------------------------------------
    //  Simple execution trace: PC + instruction
    // -------------------------------------------------
    always @(posedge clk) begin
        // Only print when the core is actually running
        if (dut.enable_design) begin
            $display("[%0t] CYCLE=%0d  PC=%08h  INSTR=%08h",
                     $time,
                     dut.Cycle_count,
                     dut.u_riscv32i_main.pc.PC,
                     dut.u_riscv32i_main.instruction);
        end
    end



    // -----------------------------------------
    // STOP_sim handling
    // -----------------------------------------
//    always @(posedge STOP_sim) begin
 //       $display("STOP_sim asserted: SUCCESS");
  //      $finish;
    //end

    // -------------------------------------------------
    //  STOP_sim handling
    // -------------------------------------------------
    always @(posedge STOP_sim) begin
        $display("STOP_sim asserted : SUCCESS");
        $display("  Cycle_count   = %0d", dut.Cycle_count);
        $display("  success_code  = 0x%08h", dut.success_code);
        $display("  final_value   = 0x%08h",
                 dut.u_riscv32i_main.dataMem.final_value);
        $finish;
    end


    always @(posedge clk) begin
        if (dut.enable_design) begin
            $display("  x1=%08h  x2=%08h  x10=%08h",
                     dut.u_riscv32i_main.reg_file.REG_FILE[1],
                     dut.u_riscv32i_main.reg_file.REG_FILE[2],
                     dut.u_riscv32i_main.reg_file.REG_FILE[10]);
        end
    end

always @(dut.u_riscv32i_main.final_value) begin
    $display("FINAL_VALUE CHANGE: %h at time %t",
             dut.u_riscv32i_main.final_value, $time);
end


    // -----------------------------------------
    // BRAM instances
    // -----------------------------------------
    bram_mem #(.MEM_DEPTH(4096)) data_mem_bram (
        .clkb(data_mem_clkb),
        .addrb(data_mem_addrb),
        .dinb(data_mem_dinb),
        .enb(data_mem_enb),
        .rstb(data_mem_rstb),
        .web(data_mem_web),
        .doutb(data_mem_doutb),
        .rstb_busy(data_mem_rstb_busy)
    );

    bram_ins #(.MEM_DEPTH(2048)) ins_mem_bram (
        .clkb(ins_mem_clkb),
        .addrb(ins_mem_addrb),
        .dinb(ins_mem_dinb),
        .enb(ins_mem_enb),
        .rstb(ins_mem_rstb),
        .web(ins_mem_web),
        .doutb(ins_mem_doutb),
        .rstb_busy(ins_mem_rstb_busy)
    );

endmodule


// =============================================================
// Data Memory BRAM
// =============================================================
module bram_mem #(parameter MEM_DEPTH = 4096) (
    input  wire        clkb,
    input  wire        enb,
    input  wire        rstb,
    input  wire [3:0]  web,
    input  wire [31:0] addrb,
    input  wire [31:0] dinb,
    output wire        rstb_busy,
    output reg [31:0]  doutb
);

    reg [31:0] DMEM [0:MEM_DEPTH-1];
    integer i;

    assign rstb_busy = 1'b0;

    initial begin
        for (i = 0; i < MEM_DEPTH; i++)
            DMEM[i] = 32'h0;
    end

    always @(posedge clkb) begin
        if (rstb) begin
            for (i = 0; i < MEM_DEPTH; i++)
                DMEM[i] <= 32'h0;
            doutb <= 32'h0;
        end else if (enb) begin
            if (web != 4'b0000) begin
                if (web[0]) DMEM[addrb[31:2]][ 7: 0] <= dinb[ 7: 0];
                if (web[1]) DMEM[addrb[31:2]][15: 8] <= dinb[15: 8];
                if (web[2]) DMEM[addrb[31:2]][23:16] <= dinb[23:16];
                if (web[3]) DMEM[addrb[31:2]][31:24] <= dinb[31:24];
            end
            doutb <= DMEM[addrb[31:2]];
        end
    end
endmodule


// =============================================================
// Instruction Memory BRAM
// =============================================================
module bram_ins #(parameter MEM_DEPTH = 2048) (
    input  wire        clkb,
    input  wire        enb,
    input  wire        rstb,
    input  wire [3:0]  web,
    input  wire [31:0] addrb,
    input  wire [31:0] dinb,
    output wire        rstb_busy,
    output reg [31:0]  doutb
);

    reg [31:0] DMEM [0:MEM_DEPTH-1];
    integer i;

    assign rstb_busy = 1'b0;

    initial begin
        for (i = 0; i < MEM_DEPTH; i++)
            DMEM[i] = 32'h00000013;

        $display("Loading program.hex into instruction memory...");
        $readmemh("program.hex", DMEM);
    end

    always @(posedge clkb) begin
        if (rstb) begin
            doutb <= 32'h0;
        end else if (enb) begin
            if (web != 4'b0000) begin
                if (web[0]) DMEM[addrb[31:2]][ 7: 0] <= dinb[ 7: 0];
                if (web[1]) DMEM[addrb[31:2]][15: 8] <= dinb[15: 8];
                if (web[2]) DMEM[addrb[31:2]][23:16] <= dinb[23:16];
                if (web[3]) DMEM[addrb[31:2]][31:24] <= dinb[31:24];
            end
            doutb <= DMEM[addrb[31:2]];
        end
    end
endmodule

