module dec_swc_wrapper (
    input hclk,
    input hrstn,
    input [3:0] cycle_cnt,
    input ifu_dec_stall,
    input [31:0] inst_in,
    output reg [31:0] inst_out,
    output reg dec_lui,
    output reg dec_auipc,
    output reg dec_jal,
    output reg dec_jalr,
    output reg dec_beq,
    output reg dec_bne,
    output reg dec_blt,
    output reg dec_bge,
    output reg dec_bltu,
    output reg dec_bgeu,
    output reg dec_lb,
    output reg dec_lh,
    output reg dec_lw,
    output reg dec_lbu,
    output reg dec_lhu,
    output reg dec_sb,
    output reg dec_sh,
    output reg dec_sw,
    output reg dec_addi,
    output reg dec_slti,
    output reg dec_sltiu,
    output reg dec_xori,
    output reg dec_ori,
    output reg dec_andi,
    output reg dec_slli,
    output reg dec_srli,
    output reg dec_srai,
    output reg dec_add,
    output reg dec_sub,
    output reg dec_sll,
    output reg dec_slt,
    output reg dec_sltu,
    output reg dec_xor,
    output reg dec_srl,
    output reg dec_sra,
    output reg dec_or,
    output reg dec_and,
    output reg dec_fence,
    output reg dec_fence_i,
    output reg dec_ecall,
    output reg dec_ebreak,
    output reg dec_csrrw,
    output reg dec_csrrs,
    output reg dec_csrrc,
    output reg dec_csrrwi,
    output reg dec_csrrsi,
    output reg dec_csrrci,
    output reg dec_upper_en,
    output reg dec_imm_en,
    output reg dec_reg_en,
    output reg dec_jump_en,
    output reg dec_branch_en,
    output reg dec_load_en,
    output reg dec_store_en,
    output reg [4:0] dec_rs2,
    output reg [4:0] dec_rs1,
    output reg [4:0] dec_rd,
    output reg [11:0] dec_imm_type_i,
    output reg [11:0] dec_imm_type_s,
    output reg [12:0] dec_imm_type_b,
    output reg [19:0] dec_imm_type_u,
    output reg [20:0] dec_imm_type_j
);

    dec_swc dut (
        .hclk(hclk),
        .hrstn(hrstn),
        .cycle_cnt(cycle_cnt),
        .ifu_dec_stall(ifu_dec_stall),
        .inst_in(inst_in),
        .inst_out(inst_out),
        .dec_lui(dec_lui),
        .dec_auipc(dec_auipc),
        .dec_jal(dec_jal),
        .dec_jalr(dec_jalr),
        .dec_beq(dec_beq),
        .dec_bne(dec_bne),
        .dec_blt(dec_blt),
        .dec_bge(dec_bge),
        .dec_bltu(dec_bltu),
        .dec_bgeu(dec_bgeu),
        .dec_lb(dec_lb),
        .dec_lh(dec_lh),
        .dec_lw(dec_lw),
        .dec_lbu(dec_lbu),
        .dec_lhu(dec_lhu),
        .dec_sb(dec_sb),
        .dec_sh(dec_sh),
        .dec_sw(dec_sw),
        .dec_addi(dec_addi),
        .dec_slti(dec_slti),
        .dec_sltiu(dec_sltiu),
        .dec_xori(dec_xori),
        .dec_ori(dec_ori),
        .dec_andi(dec_andi),
        .dec_slli(dec_slli),
        .dec_srli(dec_srli),
        .dec_srai(dec_srai),
        .dec_add(dec_add),
        .dec_sub(dec_sub),
        .dec_sll(dec_sll),
        .dec_slt(dec_slt),
        .dec_sltu(dec_sltu),
        .dec_xor(dec_xor),
        .dec_srl(dec_srl),
        .dec_sra(dec_sra),
        .dec_or(dec_or),
        .dec_and(dec_and),
        .dec_fence(dec_fence),
        .dec_fence_i(dec_fence_i),
        .dec_ecall(dec_ecall),
        .dec_ebreak(dec_ebreak),
        .dec_csrrw(dec_csrrw),
        .dec_csrrs(dec_csrrs),
        .dec_csrrc(dec_csrrc),
        .dec_csrrwi(dec_csrrwi),
        .dec_csrrsi(dec_csrrsi),
        .dec_csrrci(dec_csrrci),
        .dec_upper_en(dec_upper_en),
        .dec_imm_en(dec_imm_en),
        .dec_reg_en(dec_reg_en),
        .dec_jump_en(dec_jump_en),
        .dec_branch_en(dec_branch_en),
        .dec_load_en(dec_load_en),
        .dec_store_en(dec_store_en),
        .dec_rs2(dec_rs2),
        .dec_rs1(dec_rs1),
        .dec_rd(dec_rd),
        .dec_imm_type_i(dec_imm_type_i),
        .dec_imm_type_s(dec_imm_type_s),
        .dec_imm_type_b(dec_imm_type_b),
        .dec_imm_type_u(dec_imm_type_u),
        .dec_imm_type_j(dec_imm_type_j)
    );
    
endmodule
