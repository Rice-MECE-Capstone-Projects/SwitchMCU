// exec_driver.sv
`timescale 1ns/1ps
 import uvm_pkg::*;
import pkg_tx::*; 
`include "uvm_macros.svh"
`include "params.sv"
//`include "pkg_tx.sv"

class exec_driver extends uvm_driver #(pkg_tx::exec_tx);
  `uvm_component_utils(exec_driver)

  // virtual interface
  virtual execute_if vif;

  // publish expected transactions to scoreboard
  uvm_analysis_port#(pkg_tx::exec_tx) expected_ap;

  function new(string name, uvm_component parent);
    super.new(name, parent);
    expected_ap = new("expected_ap", this);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    // get the virtual interface (must be set from the TB)
    if (!uvm_config_db#(virtual execute_if)::get(this, "", "vif", vif)) begin
      `uvm_error("DRV", "virtual interface not found in config_db")
    end
  endfunction

  task run_phase(uvm_phase phase);
    pkg_tx::exec_tx req;
    logic [31:0] g1, g2;
      bit gb, gj, gw;
    forever begin
      // get next sequence item
      seq_item_port.get_next_item(req);
      // drive DUT pins (we assume DUT reacts combinationally, so we wait a little)
      vif.i_en = req.i_en;
      vif.rd_i = req.rd_i;
      vif.rs1_i = req.rs1_i;
      vif.rs2_i = req.rs2_i;
      vif.instruction = req.instruction;
      vif.operand1_pi = req.operand1_pi;
      vif.operand2_pi = req.operand2_pi;
      vif.imm_i = req.imm_i;
      vif.pc_i = req.pc_i;
      vif.Noop = req.Noop;
      vif.Single_Instruction_i = req.Single_Instruction_i;

      // small settling time (combinational DUT)
      @(posedge vif.clk);
      #1;

      // compute expected with golden model
      
      golden_execute(req, g1, g2, gb, gj, gw);
      req.expected_alu1 = g1;
      req.expected_alu2 = g2;
      req.expected_branch = gb;
      req.expected_jump = gj;
      req.expected_write = gw;
      req.is_expected = 1;

      // publish expected to scoreboard
      expected_ap.write(req);

      // finish the item
      seq_item_port.item_done();
    end
  endtask
endclass : exec_driver
