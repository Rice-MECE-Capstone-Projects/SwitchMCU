// pc_test.sv
`include "uvm_macros.svh"
import uvm_pkg::*;
`include "pc_env.sv"
`include "pc_seq.sv"

class pc_test extends uvm_test;
  `uvm_component_utils(pc_test)

  pc_env env;

  function new(string name="pc_test", uvm_component parent=null);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    env = pc_env::type_id::create("env", this);
  endfunction

  task run_phase(uvm_phase phase);
    pc_seq seq;
    seq = pc_seq::type_id::create("seq");
    phase.raise_objection(this);
    seq.start(env.seqr);
    #1000;  // run for 100 time units
    phase.drop_objection(this);
  endtask
endclass

