// Code your testbench here
// or browse Examples
//HELLO

`timescale 1ns/1ps
`include "params.sv" // if you need the inst_* macros
module tb_top;
  // clock
  bit clk = 0;
  always #5 clk = ~clk;

  // instantiate interface
  execute_if dut_if(.clk(clk));

  // instantiate DUT and connect to the interface signals
  execute dut0 (
    //.i_clk(clk),
    .i_en(dut_if.i_en),
    .rd_i(dut_if.rd_i),
    .rs1_i(dut_if.rs1_i),
    .rs2_i(dut_if.rs2_i),
    .instruction(dut_if.instruction),
    .operand1_pi(dut_if.operand1_pi),
    .operand2_pi(dut_if.operand2_pi),
    .imm_i(dut_if.imm_i),
    .pc_i(dut_if.pc_i),
    .Noop(dut_if.Noop),
    .alu_result_1(dut_if.alu_result_1),
    .alu_result_2(dut_if.alu_result_2),
    .branch_inst_wire(dut_if.branch_inst_wire),
    .jump_inst_wire(dut_if.jump_inst_wire),
    .write_reg_file_wire(dut_if.write_reg_file_wire),
    .Single_Instruction_i(dut_if.Single_Instruction_i)
  );

  initial begin
    // small directed smoke test
    dut_if.i_en = 1;
    dut_if.operand1_pi = 32'd10;
    dut_if.operand2_pi = 32'd7;
    dut_if.pc_i = 32'h1000;
    dut_if.imm_i = 32'd0;
    dut_if.Single_Instruction_i = `inst_ADD;
    #10;
    $display("SMOKE: alu1=%0d alu2=%0d br=%b jump=%b wr=%b", dut_if.alu_result_1, dut_if.alu_result_2, dut_if.branch_inst_wire, dut_if.jump_inst_wire, dut_if.write_reg_file_wire);
    #20 $finish;
  end
endmodule

