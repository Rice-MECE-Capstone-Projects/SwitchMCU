module top_module (
    input input hclk,
    input input hrstn,
    input input [3:0] cycle_cnt,
    input input hready,
    input input hresp,
    input input [31:0] hrdata,
    input input [4:0] exu_load_rd,
    input input [31:0] exu_load_base_addr,
    input input [31:0] exu_load_offset,
    input input exu_load_sext,
    input input [1:0] exu_load_size,
    input input exu_load_en,
    input input [31:0] exu_store_addr,
    input input [31:0] exu_store_data,
    input input exu_store_en,
    input input [1:0] exu_store_size,
    input input hclk,
    input input hrstn,
    input input hready,
    input input hresp,
    input input [31:0] hrdata,
    input input itcm_ready,
    input input ifu_dec_stall,
    input input reg [3:0] cycle_cnt,
    input input pc_write,
    input input [31:0] pc_wdata,

    output reg [31:0] haddr,
    output reg hwrite,
    output reg [31:0] hwdata,
    output reg [2:0] hsize,
    output reg [2:0] hburst,
    output reg [6:0] hprot,
    output reg [1:0] htrans,
    output reg hmastlock,
    output reg [4:0] mau_load_rd,
    output reg [31:0] mau_load_data,
    output reg mau_load_en,
    output reg [31:0] haddr,
    output hwrite,
    output reg [31:0] hwdata,
    output reg [2:0] hsize,
    output reg [2:0] hburst,
    output reg [6:0] hprot,
    output reg [1:0] htrans,
    output reg hmastlock,
    output reg ifu_idle,
    output reg [31:0] pc,
    output reg [31:0] inst_out
);


    mau_swc mau_swc_inst (
        .hclk(hclk),
        .hrstn(hrstn),
        .cycle_cnt(cycle_cnt),
        .hready(hready),
        .hresp(hresp),
        .hrdata(hrdata),
        .exu_load_rd(exu_load_rd),
        .exu_load_base_addr(exu_load_base_addr),
        .exu_load_offset(exu_load_offset),
        .exu_load_sext(exu_load_sext),
        .exu_load_size(exu_load_size),
        .exu_load_en(exu_load_en),
        .exu_store_addr(exu_store_addr),
        .exu_store_data(exu_store_data),
        .exu_store_en(exu_store_en),
        .exu_store_size(exu_store_size),
        .haddr(haddr),
        .hwrite(hwrite),
        .hwdata(hwdata),
        .hsize(hsize),
        .hburst(hburst),
        .hprot(hprot),
        .htrans(htrans),
        .hmastlock(hmastlock),
        .mau_load_rd(mau_load_rd),
        .mau_load_data(mau_load_data),
        .mau_load_en(mau_load_en)
    );

    ifu_swc ifu_swc_inst (
        .hclk(hclk),
        .hrstn(hrstn),
        .hready(hready),
        .hresp(hresp),
        .hrdata(hrdata),
        .itcm_ready(itcm_ready),
        .ifu_dec_stall(ifu_dec_stall),
        .cycle_cnt(cycle_cnt),
        .pc_write(pc_write),
        .pc_wdata(pc_wdata),
        .haddr(haddr),
        .hwrite(hwrite),
        .hwdata(hwdata),
        .hsize(hsize),
        .hburst(hburst),
        .hprot(hprot),
        .htrans(htrans),
        .hmastlock(hmastlock),
        .ifu_idle(ifu_idle),
        .pc(pc),
        .inst_out(inst_out)
    );

    initial begin
        $dumpfile("./vcds/top_module.vcd");
        $dumpvars(0, top_module);
    end
endmodule
