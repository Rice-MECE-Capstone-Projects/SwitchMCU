package core_smoke_test_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "core_smoke_test.sv"

endpackage

