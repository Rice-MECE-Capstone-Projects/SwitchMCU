module top_module (
    input input hclk,
    input input hrstn,
    input input [31:0] inst_in,
    input input dec_lui,
    input input dec_auipc,
    input input dec_jal,
    input input dec_jalr,
    input input dec_beq,
    input input dec_bne,
    input input dec_blt,
    input input dec_bge,
    input input dec_bltu,
    input input dec_bgeu,
    input input dec_lb,
    input input dec_lh,
    input input dec_lw,
    input input dec_lbu,
    input input dec_lhu,
    input input dec_sb,
    input input dec_sh,
    input input dec_sw,
    input input dec_addi,
    input input dec_slti,
    input input dec_sltiu,
    input input dec_xori,
    input input dec_ori,
    input input dec_andi,
    input input dec_slli,
    input input dec_srli,
    input input dec_srai,
    input input dec_add,
    input input dec_sub,
    input input dec_sll,
    input input dec_slt,
    input input dec_sltu,
    input input dec_xor,
    input input dec_srl,
    input input dec_sra,
    input input dec_or,
    input input dec_and,
    input input dec_fence,
    input input dec_fence_i,
    input input dec_ecall,
    input input dec_ebreak,
    input input dec_csrrw,
    input input dec_csrrs,
    input input dec_csrrc,
    input input dec_csrrwi,
    input input dec_csrrsi,
    input input dec_csrrci,
    input input dec_upper_en,
    input input dec_imm_en,
    input input dec_reg_en,
    input input dec_jump_en,
    input input dec_branch_en,
    input input dec_load_en,
    input input dec_store_en,
    input input [4:0] dec_rs2,
    input input [4:0] dec_rs1,
    input input [4:0] dec_rd,
    input input [11:0] dec_imm_type_i,
    input input [11:0] dec_imm_type_s,
    input input [12:0] dec_imm_type_b,
    input input [19:0] dec_imm_type_u,
    input input [20:0] dec_imm_type_j,
    input input [31:0] pc,
    input input [31:0] reg_rdata_1,
    input input [3:0] cycle_cnt,
    input input hclk,
    input input hrstn,
    input input [3:0] cycle_cnt,
    input input dec_upper_en,
    input input dec_lui,
    input input dec_auipc,
    input input [19:0] dec_imm_type_u,
    input input [4:0] dec_rd,
    input input [31:0] pc,
    input input exu_stall,
    input input hclk,
    input input hrstn,
    input input [3:0] cycle_cnt,
    input input dec_store_en,
    input input dec_sb,
    input input dec_sh,
    input input dec_sw,
    input input [11:0] dec_imm_type_s,
    input input [4:0] dec_rs1,
    input input [4:0] dec_rs2,
    input input [31:0] reg_rdata_1,
    input input [31:0] reg_rdata_2,
    input input exu_stall,
    input input hclk,
    input input hrstn,
    input input [3:0] cycle_cnt,
    input input en,
    input input dec_add,
    input input dec_sub,
    input input dec_sll,
    input input dec_slt,
    input input dec_sltu,
    input input dec_xor,
    input input dec_srl,
    input input dec_sra,
    input input dec_or,
    input input dec_and,
    input input [4:0] dec_rs1,
    input input [4:0] dec_rs2,
    input input [4:0] dec_rd,
    input input [31:0] pc,
    input input [31:0] reg_rdata_1,
    input input [31:0] reg_rdata_2,
    input input exu_stall,
    input input hclk,
    input input hrstn,
    input input [3:0] cycle_cnt,
    input input dec_load_en,
    input input dec_lb,
    input input dec_lh,
    input input dec_lw,
    input input dec_lbu,
    input input dec_lhu,
    input input [11:0] dec_imm_type_i,
    input input [4:0] dec_rd,
    input input [4:0] dec_rs1,
    input input [31:0] reg_rdata_1,
    input input hclk,
    input input hrstn,
    input input [3:0] cycle_cnt,
    input input dec_jump_en,
    input input dec_jal,
    input input dec_jalr,
    input input [11:0] dec_imm_type_i,
    input input [20:0] dec_imm_type_j,
    input input [4:0] dec_rd,
    input input [4:0] dec_rs1,
    input input [31:0] pc,
    input input [31:0] reg_rdata_1,
    input input hclk,
    input input hrstn,
    input input [3:0] cycle_cnt,
    input input dec_branch_en,
    input input dec_addi,
    input input dec_slti,
    input input dec_sltiu,
    input input dec_xori,
    input input dec_ori,
    input input dec_andi,
    input input dec_slli,
    input input dec_srli,
    input input dec_srai,
    input input [11:0] dec_imm_type_i,
    input input [4:0] dec_rd,
    input input [4:0] dec_rs1,
    input input [31:0] pc,
    input input [31:0] reg_rdata_1,
    input input hclk,
    input input hrstn,
    input input [3:0] cycle_cnt,
    input input [1:0] flush,
    input input hclk,
    input input hrstn,
    input input [3:0] cycle_cnt,
    input input dec_branch_en,
    input input dec_beq,
    input input dec_bne,
    input input dec_blt,
    input input dec_bge,
    input input dec_bltu,
    input input dec_bgeu,
    input input [11:0] dec_imm_type_b,
    input input [4:0] dec_rs1,
    input input [4:0] dec_rs2,
    input input [31:0] pc,
    input input [31:0] reg_rdata_1,
    input input [31:0] reg_rdata_2,

    output reg [31:0] inst_out,
    output pc_write,
    output [31:0] pc_wdata,
    output [4:0] exu_load_rd,
    output [31:0] exu_load_base_addr,
    output [31:0] exu_load_offset,
    output exu_load_sext,
    output [1:0] exu_load_size,
    output exu_load_en,
    output [31:0] exu_store_addr,
    output [31:0] exu_store_data,
    output [1:0] exu_store_size,
    output exu_store_en,
    output [4:0] reg_waddr,
    output [31:0] reg_wdata,
    output reg_wen,
    output [4:0] reg_raddr_1,
    output reg_ren_1,
    output [4:0] reg_raddr_2,
    output [31:0] reg_rdata_2,
    output reg_ren_2,
    output ifu_dec_stall,
    output reg [31:0] exu_store_addr,
    output reg [31:0] exu_store_data,
    output reg exu_store_en,
    output reg [1:0] exu_store_size,
    output ifu_dec_stall,
    output reg [4:0] exu_load_rd,
    output reg [31:0] exu_load_base_addr,
    output reg [31:0] exu_load_offset,
    output reg exu_load_sext,
    output reg [1:0] exu_load_size,
    output reg exu_load_en,
    output reg flush_stall
);


    exu_top_swc exu_top_swc_inst (
        .hclk(hclk),
        .hrstn(hrstn),
        .inst_in(inst_in),
        .dec_lui(dec_lui),
        .dec_auipc(dec_auipc),
        .dec_jal(dec_jal),
        .dec_jalr(dec_jalr),
        .dec_beq(dec_beq),
        .dec_bne(dec_bne),
        .dec_blt(dec_blt),
        .dec_bge(dec_bge),
        .dec_bltu(dec_bltu),
        .dec_bgeu(dec_bgeu),
        .dec_lb(dec_lb),
        .dec_lh(dec_lh),
        .dec_lw(dec_lw),
        .dec_lbu(dec_lbu),
        .dec_lhu(dec_lhu),
        .dec_sb(dec_sb),
        .dec_sh(dec_sh),
        .dec_sw(dec_sw),
        .dec_addi(dec_addi),
        .dec_slti(dec_slti),
        .dec_sltiu(dec_sltiu),
        .dec_xori(dec_xori),
        .dec_ori(dec_ori),
        .dec_andi(dec_andi),
        .dec_slli(dec_slli),
        .dec_srli(dec_srli),
        .dec_srai(dec_srai),
        .dec_add(dec_add),
        .dec_sub(dec_sub),
        .dec_sll(dec_sll),
        .dec_slt(dec_slt),
        .dec_sltu(dec_sltu),
        .dec_xor(dec_xor),
        .dec_srl(dec_srl),
        .dec_sra(dec_sra),
        .dec_or(dec_or),
        .dec_and(dec_and),
        .dec_fence(dec_fence),
        .dec_fence_i(dec_fence_i),
        .dec_ecall(dec_ecall),
        .dec_ebreak(dec_ebreak),
        .dec_csrrw(dec_csrrw),
        .dec_csrrs(dec_csrrs),
        .dec_csrrc(dec_csrrc),
        .dec_csrrwi(dec_csrrwi),
        .dec_csrrsi(dec_csrrsi),
        .dec_csrrci(dec_csrrci),
        .dec_upper_en(dec_upper_en),
        .dec_imm_en(dec_imm_en),
        .dec_reg_en(dec_reg_en),
        .dec_jump_en(dec_jump_en),
        .dec_branch_en(dec_branch_en),
        .dec_load_en(dec_load_en),
        .dec_store_en(dec_store_en),
        .dec_rs2(dec_rs2),
        .dec_rs1(dec_rs1),
        .dec_rd(dec_rd),
        .dec_imm_type_i(dec_imm_type_i),
        .dec_imm_type_s(dec_imm_type_s),
        .dec_imm_type_b(dec_imm_type_b),
        .dec_imm_type_u(dec_imm_type_u),
        .dec_imm_type_j(dec_imm_type_j),
        .pc(pc),
        .reg_rdata_1(reg_rdata_1),
        .cycle_cnt(cycle_cnt),
        .inst_out(inst_out),
        .pc_write(pc_write),
        .pc_wdata(pc_wdata),
        .exu_load_rd(exu_load_rd),
        .exu_load_base_addr(exu_load_base_addr),
        .exu_load_offset(exu_load_offset),
        .exu_load_sext(exu_load_sext),
        .exu_load_size(exu_load_size),
        .exu_load_en(exu_load_en),
        .exu_store_addr(exu_store_addr),
        .exu_store_data(exu_store_data),
        .exu_store_size(exu_store_size),
        .exu_store_en(exu_store_en),
        .reg_waddr(reg_waddr),
        .reg_wdata(reg_wdata),
        .reg_wen(reg_wen),
        .reg_raddr_1(reg_raddr_1),
        .reg_ren_1(reg_ren_1),
        .reg_raddr_2(reg_raddr_2),
        .reg_rdata_2(reg_rdata_2),
        .reg_ren_2(reg_ren_2),
        .ifu_dec_stall(ifu_dec_stall)
    );

    exu_upper_swc exu_upper_swc_inst (
        .hclk(hclk),
        .hrstn(hrstn),
        .cycle_cnt(cycle_cnt),
        .dec_upper_en(dec_upper_en),
        .dec_lui(dec_lui),
        .dec_auipc(dec_auipc),
        .dec_imm_type_u(dec_imm_type_u),
        .dec_rd(dec_rd),
        .pc(pc),
        .exu_stall(exu_stall),
    );

    exu_store_swc exu_store_swc_inst (
        .hclk(hclk),
        .hrstn(hrstn),
        .cycle_cnt(cycle_cnt),
        .dec_store_en(dec_store_en),
        .dec_sb(dec_sb),
        .dec_sh(dec_sh),
        .dec_sw(dec_sw),
        .dec_imm_type_s(dec_imm_type_s),
        .dec_rs1(dec_rs1),
        .dec_rs2(dec_rs2),
        .reg_rdata_1(reg_rdata_1),
        .reg_rdata_2(reg_rdata_2),
        .exu_stall(exu_stall),
        .exu_store_addr(exu_store_addr),
        .exu_store_data(exu_store_data),
        .exu_store_en(exu_store_en),
        .exu_store_size(exu_store_size)
    );

    exu_reg_swc exu_reg_swc_inst (
        .hclk(hclk),
        .hrstn(hrstn),
        .cycle_cnt(cycle_cnt),
        .en(en),
        .dec_add(dec_add),
        .dec_sub(dec_sub),
        .dec_sll(dec_sll),
        .dec_slt(dec_slt),
        .dec_sltu(dec_sltu),
        .dec_xor(dec_xor),
        .dec_srl(dec_srl),
        .dec_sra(dec_sra),
        .dec_or(dec_or),
        .dec_and(dec_and),
        .dec_rs1(dec_rs1),
        .dec_rs2(dec_rs2),
        .dec_rd(dec_rd),
        .pc(pc),
        .reg_rdata_1(reg_rdata_1),
        .reg_rdata_2(reg_rdata_2),
        .exu_stall(exu_stall),
    );

    exu_load_swc exu_load_swc_inst (
        .hclk(hclk),
        .hrstn(hrstn),
        .cycle_cnt(cycle_cnt),
        .dec_load_en(dec_load_en),
        .dec_lb(dec_lb),
        .dec_lh(dec_lh),
        .dec_lw(dec_lw),
        .dec_lbu(dec_lbu),
        .dec_lhu(dec_lhu),
        .dec_imm_type_i(dec_imm_type_i),
        .dec_rd(dec_rd),
        .dec_rs1(dec_rs1),
        .reg_rdata_1(reg_rdata_1),
        .ifu_dec_stall(ifu_dec_stall),
        .exu_load_rd(exu_load_rd),
        .exu_load_base_addr(exu_load_base_addr),
        .exu_load_offset(exu_load_offset),
        .exu_load_sext(exu_load_sext),
        .exu_load_size(exu_load_size),
        .exu_load_en(exu_load_en)
    );

    exu_jump_swc exu_jump_swc_inst (
        .hclk(hclk),
        .hrstn(hrstn),
        .cycle_cnt(cycle_cnt),
        .dec_jump_en(dec_jump_en),
        .dec_jal(dec_jal),
        .dec_jalr(dec_jalr),
        .dec_imm_type_i(dec_imm_type_i),
        .dec_imm_type_j(dec_imm_type_j),
        .dec_rd(dec_rd),
        .dec_rs1(dec_rs1),
        .pc(pc),
        .reg_rdata_1(reg_rdata_1),
    );

    exu_imm_swc exu_imm_swc_inst (
        .hclk(hclk),
        .hrstn(hrstn),
        .cycle_cnt(cycle_cnt),
        .dec_branch_en(dec_branch_en),
        .dec_addi(dec_addi),
        .dec_slti(dec_slti),
        .dec_sltiu(dec_sltiu),
        .dec_xori(dec_xori),
        .dec_ori(dec_ori),
        .dec_andi(dec_andi),
        .dec_slli(dec_slli),
        .dec_srli(dec_srli),
        .dec_srai(dec_srai),
        .dec_imm_type_i(dec_imm_type_i),
        .dec_rd(dec_rd),
        .dec_rs1(dec_rs1),
        .pc(pc),
        .reg_rdata_1(reg_rdata_1),
    );

    exu_flush_swc exu_flush_swc_inst (
        .hclk(hclk),
        .hrstn(hrstn),
        .cycle_cnt(cycle_cnt),
        .flush(flush),
        .flush_stall(flush_stall)
    );

    exu_branch_swc exu_branch_swc_inst (
        .hclk(hclk),
        .hrstn(hrstn),
        .cycle_cnt(cycle_cnt),
        .dec_branch_en(dec_branch_en),
        .dec_beq(dec_beq),
        .dec_bne(dec_bne),
        .dec_blt(dec_blt),
        .dec_bge(dec_bge),
        .dec_bltu(dec_bltu),
        .dec_bgeu(dec_bgeu),
        .dec_imm_type_b(dec_imm_type_b),
        .dec_rs1(dec_rs1),
        .dec_rs2(dec_rs2),
        .pc(pc),
        .reg_rdata_1(reg_rdata_1),
        .reg_rdata_2(reg_rdata_2),
    );

    initial begin
        $dumpfile("./vcds/top_module.vcd");
        $dumpvars(0, top_module);
    end
endmodule
