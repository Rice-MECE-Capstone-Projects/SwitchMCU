
// pc_driver.sv
`include "uvm_macros.svh"
`include "pc_txn.sv"

import uvm_pkg::*;

class pc_driver extends uvm_driver #(pc_txn);
  virtual pc_if.drv_mp vif;  // virtual interface handle

  `uvm_component_utils(pc_driver)

  function new(string name="pc_driver", uvm_component parent=null);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    if ( !uvm_config_db#(virtual pc_if.drv_mp)::get(this, "", "vif", vif) )
      `uvm_fatal("NOVIF", "virtual interface not set for pc_driver");
  endfunction


  task run_phase(uvm_phase phase);
    pc_txn tr;
    forever begin
      // Wait for a new transaction
      seq_item_port.get_next_item(tr);

      // Drive DUT inputs
      vif.stage_IF_ready   <= tr.stage_IF_ready;
      vif.jump_inst_wire   <= tr.jump_inst_wire;
      vif.branch_inst_wire <= tr.branch_inst_wire;
      vif.branch_pred_wire <= tr.branch_pred_wire;
      vif.branch_pred_old2 <= tr.branch_pred_old2;
      vif.enable_design    <= tr.enable_design;
      vif.targetPC_i       <= tr.targetPC_i;
      vif.initial_pc_i     <= tr.initial_pc_i;

      // Hold values for one clock cycle
      @(posedge vif.clk);

      // Tell UVM we're done with this transaction
      seq_item_port.item_done();
    end
  endtask
endclass
