// env.sv
`timescale 1ns/1ps
import uvm_pkg::*;
import pkg_tx::*; 
`include "uvm_macros.svh"
//`include "pkg_tx.sv"
`include "exec_driver.sv"
`include "exec_monitor.sv"
`include "exec_scoreboard.sv"

class exec_agent extends uvm_component;
  `uvm_component_utils(exec_agent)

  uvm_sequencer#(pkg_tx::exec_tx) sequencer;
  exec_driver      driver;
  exec_monitor     monitor;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    sequencer = uvm_sequencer#(pkg_tx::exec_tx)::type_id::create("sequencer", this);
    driver    = exec_driver::type_id::create("driver", this);
    monitor   = exec_monitor::type_id::create("monitor", this);
  endfunction

  function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    driver.seq_item_port.connect(sequencer.seq_item_export);
    // connect TLMs to scoreboard in ENV (the env will connect them)
  endfunction
endclass

class exec_env extends uvm_env;
  `uvm_component_utils(exec_env)

  exec_agent     agent;
  exec_scoreboard scoreboard;

  function new(string name, uvm_component parent);
    super.new(name, parent);
  endfunction

  function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    agent = exec_agent::type_id::create("agent", this);
    scoreboard = exec_scoreboard::type_id::create("scoreboard", this);
  endfunction

  function void connect_phase(uvm_phase phase);
    super.connect_phase(phase);
    // connect driver's expected port to scoreboard expected_imp
    agent.driver.expected_ap.connect(scoreboard.expected_imp);
    // connect monitor's observed port to scoreboard observed_imp
    agent.monitor.observed_ap.connect(scoreboard.observed_imp);
  endfunction
endclass
