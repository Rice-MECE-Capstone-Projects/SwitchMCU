// pc_pkg.sv
package pc_pkg;

  // Pull in UVM
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  // Include all class files here
  `include "pc_txn.sv"
  `include "pc_driver.sv"
  // later we will add:
  // `include "pc_seq.sv"
  // `include "pc_env.sv"
  // `include "pc_test.sv"

endpackage